module main;

    reg [63:0] y0;
    reg [63:0] y1;
    reg [63:0] y2;
    reg [63:0] y3;
    reg [1:0] x;
    wire [63:0] z;

    uut mux64_4_2(
        .y0(y0),
        .y1(y1),
        .y2(y2),
        .y3(y3),
        .x(x),
        .z(z)
    );

    initial begin
        // Тест 1: x = 2'b00 (y0 должно быть выбрано)
        y0 = 64'b1010101010101010101010101010101010101010101010101010101010101010;
        y1 = 64'b0101010101010101010101010101010101010101010101010101010101010101;
        y2 = 64'b1100110011001100110011001100110011001100110011001100110011001100;
        y3 = 64'b0011001100110011001100110011001100110011001100110011001100110011;
        x = 2'b00;
        #10;

        // Тест 2: x = 2'b01 (y1 должно быть выбрано)
        y0 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        y1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        y2 = 64'b1010101010101010101010101010101010101010101010101010101010101010;
        y3 = 64'b0101010101010101010101010101010101010101010101010101010101010101;
        x = 2'b01;
        #10;

        // Тест 3: x = 2'b10 (y2 должно быть выбрано)
        y0 = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        y1 = 64'b0100000000000000000000000000000000000000000000000000000000000000;
        y2 = 64'b0011111111111111111111111111111111111111111111111111111111111111;
        y3 = 64'b0001111111111111111111111111111111111111111111111111111111111111;
		x = 2'b10;
		#10;
      
      	// Тест 4: x = 2'b11 (y3 должно быть выбрано)
        y0 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        y1 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        y2 = 64'b1111000011110000111100001111000011110000111100001111000011110000;
        y3 = 64'b0000111100001111000011110000111100001111000011110000111100001111;
        x = 2'b11;
        #10;

      end;
endmodule


